function Bit#(8) charToAscii(Char c);
  case (c) matches
    "0" : return 48;
    "1" : return 49;
    "2" : return 50;
    "3" : return 51;
    "4" : return 52;
    "5" : return 53;
    "6" : return 54;
    "7" : return 55;
    "8" : return 56;
    "9" : return 57;
    "a" : return 97;
    "b" : return 98;
    "c" : return 99;
    "d" : return 100;
    "e" : return 101;
    "f" : return 102;
    "g" : return 103;
    "h" : return 104;
    "i" : return 105;
    "j" : return 106;
    "k" : return 107;
    "l" : return 108;
    "m" : return 109;
    "n" : return 110;
    "o" : return 111;
    "p" : return 112;
    "q" : return 113;
    "r" : return 114;
    "s" : return 115;
    "t" : return 116;
    "u" : return 117;
    "v" : return 118;
    "w" : return 119;
    "x" : return 120;
    "y" : return 121;
    "z" : return 122;
    "A" : return 65;
    "B" : return 66;
    "C" : return 67;
    "D" : return 68;
    "E" : return 69;
    "F" : return 70;
    "G" : return 71;
    "H" : return 72;
    "I" : return 73;
    "J" : return 74;
    "K" : return 75;
    "L" : return 76;
    "M" : return 77;
    "N" : return 78;
    "O" : return 79;
    "P" : return 80;
    "Q" : return 81;
    "R" : return 82;
    "S" : return 83;
    "T" : return 84;
    "U" : return 85;
    "V" : return 86;
    "W" : return 87;
    "X" : return 88;
    "Y" : return 89;
    "Z" : return 90;
    "!" : return 33;
    "\"" : return 34;
    "#" : return 35;
    "$" : return 36;
    "%" : return 37;
    "&" : return 38;
    "'" : return 39;
    "(" : return 40;
    ")" : return 41;
    "*" : return 42;
    "+" : return 43;
    "," : return 44;
    "-" : return 45;
    "." : return 46;
    "/" : return 47;
    ":" : return 58;
    ";" : return 59;
    "<" : return 60;
    "=" : return 61;
    ">" : return 62;
    "?" : return 63;
    "@" : return 64;
    "[" : return 91;
    "\\" : return 92;
    "]" : return 93;
    "^" : return 94;
    "_" : return 95;
    "{" : return 123;
    "|" : return 124;
    "}" : return 125;
    "~" : return 126;
    " " : return 32;
    "\t" : return 9;
    "\n" : return 10;
    "\x0b" : return 11;
    "\x0c" : return 12;
    default : return 95;
  endcase
endfunction
