// megafunction wizard: %10GBASE-R PHY v16.0%
// GENERATION: XML
// phy.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module phy (
		input  wire         pll_ref_clk,          //        pll_ref_clk.clk
		output wire         xgmii_rx_clk,         //       xgmii_rx_clk.clk
		output wire         pll_locked,           //         pll_locked.export
		output wire         tx_ready,             //           tx_ready.export
		input  wire         xgmii_tx_clk,         //       xgmii_tx_clk.clk
		output wire         rx_ready,             //           rx_ready.export
		output wire [3:0]   rx_data_ready,        //      rx_data_ready.export
		output wire [71:0]  xgmii_rx_dc_0,        //      xgmii_rx_dc_0.data
		input  wire         rx_serial_data_0,     //   rx_serial_data_0.export
		output wire [71:0]  xgmii_rx_dc_1,        //      xgmii_rx_dc_1.data
		input  wire         rx_serial_data_1,     //   rx_serial_data_1.export
		output wire [71:0]  xgmii_rx_dc_2,        //      xgmii_rx_dc_2.data
		input  wire         rx_serial_data_2,     //   rx_serial_data_2.export
		output wire [71:0]  xgmii_rx_dc_3,        //      xgmii_rx_dc_3.data
		input  wire         rx_serial_data_3,     //   rx_serial_data_3.export
		input  wire [71:0]  xgmii_tx_dc_0,        //      xgmii_tx_dc_0.data
		output wire [0:0]   tx_serial_data_0,     //   tx_serial_data_0.export
		input  wire [71:0]  xgmii_tx_dc_1,        //      xgmii_tx_dc_1.data
		output wire [0:0]   tx_serial_data_1,     //   tx_serial_data_1.export
		input  wire [71:0]  xgmii_tx_dc_2,        //      xgmii_tx_dc_2.data
		output wire [0:0]   tx_serial_data_2,     //   tx_serial_data_2.export
		input  wire [71:0]  xgmii_tx_dc_3,        //      xgmii_tx_dc_3.data
		output wire [0:0]   tx_serial_data_3,     //   tx_serial_data_3.export
		output wire [367:0] reconfig_from_xcvr,   // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [559:0] reconfig_to_xcvr,     //   reconfig_to_xcvr.reconfig_to_xcvr
		input  wire         phy_mgmt_clk,         //       phy_mgmt_clk.clk
		input  wire         phy_mgmt_clk_reset,   // phy_mgmt_clk_reset.reset
		input  wire [8:0]   phy_mgmt_address,     //           phy_mgmt.address
		input  wire         phy_mgmt_read,        //                   .read
		output wire [31:0]  phy_mgmt_readdata,    //                   .readdata
		input  wire         phy_mgmt_write,       //                   .write
		input  wire [31:0]  phy_mgmt_writedata,   //                   .writedata
		output wire         phy_mgmt_waitrequest  //                   .waitrequest
	);

	wire    [3:0] phy_inst_tx_serial_data; // port fragment
	wire  [287:0] phy_inst_xgmii_rx_dc;    // port fragment

	altera_xcvr_10gbaser #(
		.device_family            ("Stratix V"),
		.num_channels             (4),
		.operation_mode           ("duplex"),
		.external_pma_ctrl_config (0),
		.control_pin_out          (0),
		.recovered_clk_out        (0),
		.pll_locked_out           (1),
		.ref_clk_freq             ("644.53125 MHz"),
		.pma_mode                 (40),
		.pll_type                 ("CMU"),
		.starting_channel_number  (0),
		.reconfig_interfaces      (8),
		.rx_use_coreclk           (0),
		.embedded_reset           (1),
		.latadj                   (0),
		.high_precision_latadj    (1),
		.tx_termination           ("OCT_100_OHMS"),
		.tx_vod_selection         (7),
		.tx_preemp_pretap         (0),
		.tx_preemp_pretap_inv     (0),
		.tx_preemp_tap_1          (15),
		.tx_preemp_tap_2          (0),
		.tx_preemp_tap_2_inv      (0),
		.rx_common_mode           ("0.82v"),
		.rx_termination           ("OCT_100_OHMS"),
		.rx_eq_dc_gain            (0),
		.rx_eq_ctrl               (0),
		.mgmt_clk_in_mhz          (150)
	) phy_inst (
		.pll_ref_clk          (pll_ref_clk),                                                                                                           //        pll_ref_clk.clk
		.xgmii_rx_clk         (xgmii_rx_clk),                                                                                                          //       xgmii_rx_clk.clk
		.pll_locked           (pll_locked),                                                                                                            //         pll_locked.export
		.tx_ready             (tx_ready),                                                                                                              //           tx_ready.export
		.xgmii_tx_clk         (xgmii_tx_clk),                                                                                                          //       xgmii_tx_clk.clk
		.rx_ready             (rx_ready),                                                                                                              //           rx_ready.export
		.rx_data_ready        (rx_data_ready),                                                                                                         //      rx_data_ready.export
		.xgmii_rx_dc          ({phy_inst_xgmii_rx_dc[287:216],phy_inst_xgmii_rx_dc[215:144],phy_inst_xgmii_rx_dc[143:72],phy_inst_xgmii_rx_dc[71:0]}), //      xgmii_rx_dc_0.data
		.rx_serial_data       ({rx_serial_data_3,rx_serial_data_2,rx_serial_data_1,rx_serial_data_0}),                                                 //   rx_serial_data_0.export
		.xgmii_tx_dc          ({xgmii_tx_dc_3[71:0],xgmii_tx_dc_2[71:0],xgmii_tx_dc_1[71:0],xgmii_tx_dc_0[71:0]}),                                     //      xgmii_tx_dc_0.data
		.tx_serial_data       ({phy_inst_tx_serial_data[3],phy_inst_tx_serial_data[2],phy_inst_tx_serial_data[1],phy_inst_tx_serial_data[0]}),         //   tx_serial_data_0.export
		.reconfig_from_xcvr   (reconfig_from_xcvr),                                                                                                    // reconfig_from_xcvr.reconfig_from_xcvr
		.reconfig_to_xcvr     (reconfig_to_xcvr),                                                                                                      //   reconfig_to_xcvr.reconfig_to_xcvr
		.phy_mgmt_clk         (phy_mgmt_clk),                                                                                                          //       phy_mgmt_clk.clk
		.phy_mgmt_clk_reset   (phy_mgmt_clk_reset),                                                                                                    // phy_mgmt_clk_reset.reset
		.phy_mgmt_address     (phy_mgmt_address),                                                                                                      //           phy_mgmt.address
		.phy_mgmt_read        (phy_mgmt_read),                                                                                                         //                   .read
		.phy_mgmt_readdata    (phy_mgmt_readdata),                                                                                                     //                   .readdata
		.phy_mgmt_write       (phy_mgmt_write),                                                                                                        //                   .write
		.phy_mgmt_writedata   (phy_mgmt_writedata),                                                                                                    //                   .writedata
		.phy_mgmt_waitrequest (phy_mgmt_waitrequest),                                                                                                  //                   .waitrequest
		.rx_block_lock        (),                                                                                                                      //        (terminated)
		.rx_hi_ber            (),                                                                                                                      //        (terminated)
		.rx_recovered_clk     (),                                                                                                                      //        (terminated)
		.rx_coreclkin         (1'b0),                                                                                                                  //        (terminated)
		.gxb_pdn              (1'b0),                                                                                                                  //        (terminated)
		.pll_pdn              (1'b0),                                                                                                                  //        (terminated)
		.cal_blk_pdn          (1'b0),                                                                                                                  //        (terminated)
		.cal_blk_clk          (1'b0),                                                                                                                  //        (terminated)
		.tx_digitalreset      (4'b0000),                                                                                                               //        (terminated)
		.tx_analogreset       (4'b0000),                                                                                                               //        (terminated)
		.tx_cal_busy          (),                                                                                                                      //        (terminated)
		.pll_powerdown        (4'b0000),                                                                                                               //        (terminated)
		.rx_digitalreset      (4'b0000),                                                                                                               //        (terminated)
		.rx_analogreset       (4'b0000),                                                                                                               //        (terminated)
		.rx_cal_busy          (),                                                                                                                      //        (terminated)
		.rx_is_lockedtodata   (),                                                                                                                      //        (terminated)
		.rx_latency_adj       (),                                                                                                                      //        (terminated)
		.tx_latency_adj       ()                                                                                                                       //        (terminated)
	);

	assign tx_serial_data_3 = { phy_inst_tx_serial_data[3] };

	assign xgmii_rx_dc_1 = { phy_inst_xgmii_rx_dc[143:72] };

	assign tx_serial_data_1 = { phy_inst_tx_serial_data[1] };

	assign xgmii_rx_dc_3 = { phy_inst_xgmii_rx_dc[287:216] };

	assign tx_serial_data_2 = { phy_inst_tx_serial_data[2] };

	assign xgmii_rx_dc_0 = { phy_inst_xgmii_rx_dc[71:0] };

	assign xgmii_rx_dc_2 = { phy_inst_xgmii_rx_dc[215:144] };

	assign tx_serial_data_0 = { phy_inst_tx_serial_data[0] };

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2017 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_10gbaser" version="16.0" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="num_channels" value="4" />
// Retrieval info: 	<generic name="operation_mode" value="duplex" />
// Retrieval info: 	<generic name="external_pma_ctrl_config" value="0" />
// Retrieval info: 	<generic name="control_pin_out" value="0" />
// Retrieval info: 	<generic name="recovered_clk_out" value="0" />
// Retrieval info: 	<generic name="pll_locked_out" value="1" />
// Retrieval info: 	<generic name="gui_pll_type" value="CMU" />
// Retrieval info: 	<generic name="ref_clk_freq" value="644.53125 MHz" />
// Retrieval info: 	<generic name="pma_mode" value="40" />
// Retrieval info: 	<generic name="starting_channel_number" value="0" />
// Retrieval info: 	<generic name="sys_clk_in_hz" value="150000000" />
// Retrieval info: 	<generic name="rx_use_coreclk" value="0" />
// Retrieval info: 	<generic name="gui_embedded_reset" value="1" />
// Retrieval info: 	<generic name="latadj" value="0" />
// Retrieval info: 	<generic name="high_precision_latadj" value="1" />
// Retrieval info: 	<generic name="tx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="tx_vod_selection" value="7" />
// Retrieval info: 	<generic name="tx_preemp_pretap" value="0" />
// Retrieval info: 	<generic name="tx_preemp_pretap_inv" value="0" />
// Retrieval info: 	<generic name="tx_preemp_tap_1" value="15" />
// Retrieval info: 	<generic name="tx_preemp_tap_2" value="0" />
// Retrieval info: 	<generic name="tx_preemp_tap_2_inv" value="0" />
// Retrieval info: 	<generic name="rx_common_mode" value="0.82v" />
// Retrieval info: 	<generic name="rx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="rx_eq_dc_gain" value="0" />
// Retrieval info: 	<generic name="rx_eq_ctrl" value="0" />
// Retrieval info: 	<generic name="mgmt_clk_in_hz" value="150000000" />
// Retrieval info: </instance>
// IPFS_FILES : phy.vo
// RELATED_FILES: phy.v, altera_xcvr_functions.sv, alt_reset_ctrl_lego.sv, alt_reset_ctrl_tgx_cdrauto.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_10gbaser_phy_clock_crosser.v, altera_10gbaser_phy_pipeline_stage.sv, altera_10gbaser_phy_pipeline_base.v, altera_std_synchronizer_nocut.v, csr_pcs10gbaser_h.sv, csr_pcs10gbaser.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, sv_xcvr_10gbaser_nr.sv, sv_xcvr_10gbaser_native.sv, altera_xcvr_10gbaser.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv
