`include "config.v"

// Example accelerator which consumes a message, and then sends it to the
// address specified in the first word of the message's payload.

typedef struct packed {
  logic acc;
  logic host;
  logic hostDir;
  logic [`TinselMeshYBits-1:0] boardY;
  logic [`TinselMeshXBits-1:0] boardX;
  logic [`TinselMailboxMeshYBits-1:0] tileY;
  logic [`TinselMailboxMeshXBits-1:0] tileX;
  logic [`TinselLogCoresPerMailbox-1:0] coreId;
  logic [`TinselLogThreadsPerCore-1:0] threadId;
} NetAddr;

typedef struct packed {
  // Destination address
  NetAddr dest;
  // Size of payload in 32-bit words
  logic [`TinselLogWordsPerMsg-1:0] numWords;
  // Is this a special packet for idle-detection?
  logic isIdleToken;
  // Payload
  logic [`TinselBitsPerMsg-1:0] payload;
} Msg;

module ExternalTinselAccelerator
  ( // Clock and reset
    // By default, BSV synchronises on negedge(clock) and uses negative reset
    input wire clk
  , input wire rst_n

    // Coordinates of this FPGA board in the board mesh
  , input wire [`TinselMeshXBits-1:0] board_x
  , input wire [`TinselMeshYBits-1:0] board_y

    // Stream of messages coming in
  , input wire [$bits(Msg)-1:0] in_data
  , input wire in_valid
  , output wire in_ready

    // Stream of messages going out
  , output wire [$bits(Msg)-1:0] out_data
  , output wire out_valid
  , input wire out_ready
  );

  // Compile-time NoC coordinates of this accelerator
  parameter TILE_X = 0;
  parameter TILE_Y = 0;

  // Input message queue
  reg inQueueFull = 0;
  Msg inQueueData;

  assign in_ready = !inQueueFull;

  // Output message queue
  reg outQueueFull = 0;
  Msg outQueueData;

  assign out_valid = outQueueFull;
  assign out_data = outQueueData;

  // State machine
  always @(negedge clk) begin
    if (rst_n == 0) begin
      inQueueFull <= 0;
      outQueueFull <= 0;
    end else begin
      if (in_valid && !inQueueFull) begin
        inQueueFull <= 1;
        inQueueData <= in_data;
      end

      if (outQueueFull && out_ready) begin
        outQueueFull <= 0;
      end

      if (inQueueFull && !outQueueFull) begin
        outQueueFull <= 1;
        outQueueData <= '{
            dest: inQueueData.payload[$bits(NetAddr)-1:0]
          , numWords: `TinselWordsPerMsg-1
          , isIdleToken: 0
          , payload: inQueueData.payload
        };
        inQueueFull <= 0;
      end
    end
  end

endmodule
